module bad_no_assign (
	input		a,
	input		b,
	output	y
	);
	
	wire n0;
	
//	y = ~n0;
//	n0 = a & b;
	
endmodule

