module adder4 (
	input  [3:0] a,
	input  [3:0] b,
	output [3:0] s
	);
	
	assign s = a + b;
	
endmodule
